LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.NUMERIC_STD.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY draw_map IS PORT (
    world_X, world_Y:			IN STD_LOGIC_VECTOR(8 downto 0);
    tile_num:						IN STD_LOGIC_VECTOR(2 downto 0);
    red, green, blue:			OUT STD_LOGIC
    );
END;

ARCHITECTURE bhv of draw_map IS 
	SIGNAL sub_X, sub_Y: STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL tile_addr: STD_LOGIC_VECTOR(10 downto 0);
	SIGNAL tile_data: STD_LOGIC_VECTOR(2 downto 0);
    
	SUBTYPE tile_pixel IS integer RANGE 0 TO 7;
	TYPE rom_type IS ARRAY(0 TO 2047) OF tile_pixel;
	CONSTANT tile_rom: rom_type :=
	(
		-- 0
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,

		-- 1 wood --
		6,6,6,7,0,7,0,7,7,6,6,7,7,7,6,7,
		6,6,5,6,6,0,0,0,7,7,7,6,7,7,7,6,
		6,6,5,7,7,0,6,0,0,6,6,7,7,6,7,7,
		6,6,5,7,7,6,6,6,0,0,7,7,6,7,7,6,
		7,6,5,7,7,7,6,6,6,0,0,7,6,7,7,6,
		0,6,5,7,7,7,6,5,6,6,0,0,6,6,7,6,
		0,0,7,5,7,7,6,5,7,6,6,0,0,6,7,7,
		7,0,0,5,7,7,6,6,5,6,6,6,0,0,6,6,
		7,6,0,0,7,7,6,6,5,7,7,6,0,0,0,7,
		7,0,0,0,6,7,7,6,6,5,7,0,6,6,6,0,
		7,7,6,0,0,6,7,6,6,5,0,6,7,7,7,6,
		7,7,6,0,0,0,6,7,6,0,6,7,7,6,6,6,
		7,7,6,6,5,0,0,6,7,0,6,6,6,7,6,6,
		7,7,6,6,6,5,0,0,6,0,7,7,7,7,6,6,
		7,7,7,7,6,5,7,0,0,0,6,7,7,7,7,6,
		2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,

-- 0: black
-- 1: blue 
-- 2: green
-- 3: cyan
-- 4: red
-- 5: purple
-- 6: yellow
-- 7: white
		-- 2 stone --
		3,3,3,3,3,4,3,3,4,4,3,3,3,3,3,3,
		3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,
		3,3,3,3,0,0,0,0,0,0,0,0,6,4,4,6,
		3,3,3,0,0,0,0,0,0,0,0,0,0,6,4,6,
		3,3,0,0,0,0,6,6,6,6,6,0,0,0,6,4,
		3,0,0,0,6,6,6,6,6,6,6,6,0,0,0,4,
		3,0,0,6,6,0,0,0,0,0,6,6,6,0,0,0,
		0,0,0,6,6,6,6,6,6,6,6,6,6,6,0,0,
		0,0,6,6,6,6,6,6,6,6,6,6,6,6,0,0,
		3,0,6,6,6,6,6,6,6,6,6,6,6,6,0,0,
		3,0,0,6,6,0,0,0,0,0,6,6,6,6,0,0,
		3,0,0,0,6,6,6,6,6,6,6,6,6,6,0,0,
		3,0,0,0,6,6,6,6,6,6,6,6,6,0,0,3,
		3,3,0,0,0,0,0,0,0,0,0,0,0,0,3,3,
		3,3,3,0,0,0,0,0,0,0,0,0,0,3,3,3,
		3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,


		-- 3 grass --
		0,0,0,0,0,0,0,3,0,0,0,0,0,3,0,0,
		0,0,0,0,0,0,0,2,2,0,0,0,0,2,0,0,
		0,3,0,0,0,0,0,2,2,0,0,0,0,2,0,0,
		0,2,3,0,0,0,2,2,2,2,0,0,7,3,3,2,
		0,2,3,0,0,0,2,2,2,2,0,0,3,3,2,2,
		3,2,2,0,0,3,2,2,2,2,3,0,2,3,3,2,
		3,2,2,3,0,2,2,2,2,2,2,3,2,3,4,2,
		3,2,2,2,3,2,2,2,2,2,3,2,2,2,2,2,
		3,2,2,2,3,2,2,2,2,2,3,2,2,2,2,2,
		3,2,2,2,2,2,3,2,2,2,2,2,2,2,2,2,
		2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,
		2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,
		2,2,2,2,2,2,2,2,2,3,2,2,2,2,2,2,
		2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,
		2,2,2,3,3,3,3,2,3,3,2,2,2,2,3,2,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,

		-- 4
		4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,
		4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,4,4,4,4,4,4,4,4,0,0,4,4,
		4,4,0,0,4,4,4,4,4,4,4,4,0,0,4,4,
		4,4,0,0,4,4,4,4,4,4,4,4,0,0,4,4,
		4,4,0,0,4,4,4,4,4,4,4,4,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,0,0,0,0,0,0,0,0,0,0,0,0,4,4,
		4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,
		4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,

		-- 5
		1,2,1,2,1,2,1,2,1,2,1,2,1,2,1,2,
		2,4,2,4,2,4,2,4,2,4,2,4,2,4,2,4,
		3,4,3,4,3,4,3,4,3,4,3,4,3,4,3,4,
		3,5,3,5,3,5,3,5,3,5,3,5,3,5,3,5,
		5,6,5,6,5,6,5,6,5,6,5,6,5,6,5,6,
		1,2,1,2,1,2,1,2,1,2,1,2,1,2,1,2,
		2,4,2,4,2,4,2,4,2,4,2,4,2,4,2,4,
		3,4,3,4,3,4,3,4,3,4,3,4,3,4,3,4,
		3,5,3,5,3,5,3,5,3,5,3,5,3,5,3,5,
		7,6,5,4,3,2,1,0,0,1,2,3,4,5,6,7,
		6,5,4,3,2,1,0,0,1,2,3,4,5,6,7,7,
		5,4,3,2,1,0,0,1,2,3,4,5,6,7,7,6,
		4,3,2,1,0,0,1,2,3,4,5,6,7,7,6,5,
		3,2,1,0,0,1,2,3,4,5,6,7,7,6,5,4,
		2,1,0,0,1,2,3,4,5,6,7,7,6,5,4,3,
		1,0,0,1,2,3,4,5,6,7,7,6,5,4,3,2,

		-- 6
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,4,4,4,4,0,0,0,0,0,0,
		0,0,0,0,4,4,4,4,7,4,4,4,0,0,0,0,
		0,4,4,4,4,7,7,4,4,4,4,4,4,4,4,0,
		4,4,7,4,4,7,4,4,4,7,4,4,7,4,4,4,
		4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,
		0,0,4,4,4,4,4,7,7,4,4,4,4,4,0,0,
		0,0,0,0,0,0,7,7,7,7,0,0,0,0,0,0,
		0,0,0,0,0,0,7,7,7,7,0,0,0,0,0,0,
		0,0,0,0,0,0,7,7,7,7,0,0,0,0,0,0,
		0,0,0,0,0,0,7,7,7,7,0,0,0,0,0,0,
		0,0,0,0,0,7,7,7,7,7,7,0,0,0,0,0,
		0,0,0,0,0,7,7,7,7,7,7,0,0,0,0,0,
		0,0,0,0,0,7,7,7,7,7,7,0,0,0,0,0,

		-- 7
		0,6,6,6,6,6,6,6,6,6,6,6,6,6,0,0,
		6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,0,
		6,6,1,6,6,6,0,0,0,0,6,6,1,6,6,0,
		6,6,6,6,6,0,0,6,6,0,0,6,6,6,6,0,
		6,6,6,6,0,0,6,6,6,6,0,0,6,6,6,0,
		6,6,6,6,0,0,6,6,6,6,0,0,6,6,6,0,
		6,6,6,6,6,6,6,6,6,0,0,6,6,6,6,0,
		6,6,6,6,6,6,6,6,0,0,6,6,6,6,6,0,
		6,6,6,6,6,6,6,0,0,6,6,6,6,6,6,0,
		6,6,6,6,6,6,6,0,0,6,6,6,6,6,6,0,
		6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,0,
		6,6,6,6,6,6,6,0,0,6,6,6,6,6,6,0,
		6,6,1,6,6,6,6,0,0,6,6,6,1,6,6,0,
		6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,0,
		0,6,6,6,6,6,6,6,6,6,6,6,6,6,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	);
	
	
BEGIN
	
	sub_X <= world_X(3 downto 0);
	sub_Y <= world_Y(3 downto 0);

	tile_addr <= tile_num & sub_Y & sub_X;
	
	PROCESS(tile_addr)
		VARIABLE tile: tile_pixel;
	BEGIN
	tile := tile_rom(to_integer(unsigned(tile_addr)));
	case tile is
		when 0 => tile_data <= "000";
		when 1 => tile_data <= "001";
		when 2 => tile_data <= "010";
		when 3 => tile_data <= "011";
		when 4 => tile_data <= "100";
		when 5 => tile_data <= "101";
		when 6 => tile_data <= "110";
		when 7 => tile_data <= "111";
		when others => tile_data <= "000";
	end case;
	--tile_data <= CONV_STD_LOGIC_VECTOR(, 3);
	END PROCESS;
	
	PROCESS(tile_data)
	BEGIN
		red <= tile_data(2);
		green <= tile_data(1);
		blue <= tile_data(0);
	END PROCESS;
END bhv;