LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.NUMERIC_STD.all;
--USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY map_rom IS PORT(
		clock:			IN STD_LOGIC;
		tile_X:			IN STD_LOGIC_VECTOR(4 downto 0);
		tile_Y:			IN STD_LOGIC_VECTOR(4 downto 0);
		data:				OUT STD_LOGIC_VECTOR(2 downto 0)
	);
END;

ARCHITECTURE map_rom OF map_rom IS
    SIGNAL addr: STD_LOGIC_VECTOR(9 downto 0);

    SUBTYPE map_tile IS integer RANGE 0 TO 7;
    TYPE rom_type IS ARRAY(0 TO 1023) OF map_tile;
	CONSTANT rom: rom_type :=
	(
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,7,7,7,7,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		4,4,4,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,4,4,4,0,0,0,2,0,0,0,0,0,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,2,0,0,0,0,0,0,5,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,
		0,0,0,0,0,0,0,2,0,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0,2,2,0,0,0,0,0,0,
		0,0,0,0,0,0,2,0,0,0,6,6,0,5,5,5,5,5,0,6,6,0,0,0,2,2,2,0,0,0,0,0,
		1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
		0,0,0,0,0,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0,
		0,0,0,0,0,0,0,0,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0,
		0,0,0,0,0,4,0,0,0,0,3,0,0,0,3,0,0,3,0,0,0,0,0,0,0,2,0,0,2,2,2,2,
		0,0,0,0,3,4,4,4,0,0,3,0,0,0,3,0,0,3,3,0,0,0,0,3,0,2,0,0,0,0,0,0,
		0,0,0,0,3,3,0,0,0,0,3,3,3,3,3,0,0,3,3,3,0,0,3,3,0,2,0,0,0,0,0,0,
		3,3,3,3,0,0,0,0,0,0,4,0,0,0,2,0,0,0,0,2,0,3,2,2,2,2,2,2,2,2,0,0,
		0,0,0,0,0,4,0,0,4,4,4,0,0,0,2,0,0,0,0,2,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,4,0,0,0,0,0,0,0,0,2,0,0,0,0,2,2,2,2,2,2,2,0,0,0,0,0,0,
		0,0,5,5,0,4,5,0,0,0,0,0,0,0,2,0,0,0,0,2,2,2,2,2,2,2,2,0,0,2,2,2,
		0,0,5,5,0,4,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,3,0,0,3,0,3,0,0,0,3,0,
		0,0,0,0,0,4,5,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,0,0,0,0,0,3,0,
		0,0,0,0,0,4,5,5,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,0,
		0,0,0,0,0,4,5,5,5,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,0,0,
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1
	);
BEGIN
    addr <= tile_Y & tile_X;
    
    PROCESS(clock)
		VARIABLE temp: map_tile;
    BEGIN
    	IF clock'Event AND clock = '1' THEN
			temp := rom(to_integer(unsigned(addr)));
			case temp is
				when 0 => data <= "000";
				when 1 => data <= "001";
				when 2 => data <= "010";
				when 3 => data <= "011";
				when 4 => data <= "100";
				when 5 => data <= "101";
				when 6 => data <= "110";
				when 7 => data <= "111";
				when others => data <= "000";
			end case;
	-- data <= CONV_STD_LOGIC_VECTOR(, 3);
      END IF;
    END PROCESS;
END map_rom;